`timescale 1ns / 1ps

// 32-to-5 Priority Encoder (Structural)

//behavioral model
module encoder32to5(
    input  [31:0] D,  
    output [4:0]  Y,    
    output        V   
);
    always @* begin
        V = |D;
       case (D)
           32'b0000_0000_0000_0000_0000_0000_0000_0001 : Y = 5'd0;
           32'b0000_0000_0000_0000_0000_0000_0000_0010 : Y = 5'd1;
           32'b0000_0000_0000_0000_0000_0000_0000_0100 : Y = 5'd2;
           32'b0000_0000_0000_0000_0000_0000_0000_1000 : Y = 5'd3;
           32'b0000_0000_0000_0000_0000_0000_0001_0000 : Y = 5'd4;
           32'b0000_0000_0000_0000_0000_0000_0010_0000 : Y = 5'd5;
           32'b0000_0000_0000_0000_0000_0000_0100_0000 : Y = 5'd6;
           32'b0000_0000_0000_0000_0000_0000_1000_0000 : Y = 5'd7;
           32'b0000_0000_0000_0000_0000_0001_0000_0000 : Y = 5'd8;
           32'b0000_0000_0000_0000_0000_0010_0000_0000 : Y = 5'd9;
           32'b0000_0000_0000_0000_0000_0100_0000_0000 : Y = 5'd10;
           32'b0000_0000_0000_0000_0000_1000_0000_0000 : Y = 5'd11;
           32'b0000_0000_0000_0000_0001_0000_0000_0000 : Y = 5'd12;
           32'b0000_0000_0000_0000_0010_0000_0000_0000 : Y = 5'd13;
           32'b0000_0000_0000_0000_0100_0000_0000_0000 : Y = 5'd14;
           32'b0000_0000_0000_0000_1000_0000_0000_0000 : Y = 5'd15;
           32'b0000_0000_0001_0000_0000_0000_0000_0000 : Y = 5'd16;
           32'b0000_0000_0010_0000_0000_0000_0000_0000 : Y = 5'd17;
           32'b0000_0000_0100_0000_0000_0000_0000_0000 : Y = 5'd18;
           32'b0000_0000_1000_0000_0000_0000_0000_0000 : Y = 5'd19;
           32'b0000_0001_0000_0000_0000_0000_0000_0000 : Y = 5'd20;
           32'b0000_0010_0000_0000_0000_0000_0000_0000 : Y = 5'd21;
           32'b0000_0100_0000_0000_0000_0000_0000_0000 : Y = 5'd22;
           32'b0000_1000_0000_0000_0000_0000_0000_0000 : Y = 5'd23;
           32'b0001_0000_0000_0000_0000_0000_0000_0000 : Y = 5'd24;
           32'b0010_0000_0000_0000_0000_0000_0000_0000 : Y = 5'd25;
           32'b0100_0000_0000_0000_0000_0000_0000_ 0000 : Y = 5'd26;
           32'b1000_0000_0000_0000_0000_0000_0000_0000 : Y = 5'd27;
           default: Y = 5'd0; // when none asserted or multiple asserted
       endcase
    end
endmodule
//structural model
module encoder32to5_structural (
    input  [31:0] D,  
    output [4:0]  Y,    
    output        V   
);  
    wire        v_hi, v_lo;
    wire [2:0]  y_hi, y_lo;
    
    encoder16to4_structural enc_hi (
        .D(D[31:16]),
        .Y(y_hi),
        .V(v_hi)
    );
    encoder16to4_structural enc_lo (
        .D(D[15:0]),
        .Y(y_lo),
        .V(v_lo)
    );
    assign V      = v_hi | v_lo;
    assign Y[4]   = v_hi;
    assign Y[3]   = v_hi ? y_hi[3] : y_lo[3];
    assign Y[2]   = v_hi ? y_hi[2] : y_lo[2];
    assign Y[1]   = v_hi ? y_hi[1] : y_lo[1];
    assign Y[0]   = v_hi ? y_hi[0] : y_lo[0];
endmodule

//dataflow model
module encoder32to5_dataflow (
    input  [31:0] D,  
    output [4:0]  Y,    
    output        V  
);  
    wire        v_hi, v_lo;
    wire [2:0]  y_hi, y_lo;
    
    encoder16to4_dataflow enc_hi (
        .D(D[31:16]),
        .Y(y_hi),
        .V(v_hi)
    );
    encoder16to4_dataflow enc_lo (
        .D(D[15:0]),
        .Y(y_lo),
        .V(v_lo)
    );
    assign V      = v_hi | v_lo;
    assign Y[4]   = v_hi;
    assign Y[3]   = v_hi ? y_hi[3] : y_lo[3];
    assign Y[2]   = v_hi ? y_hi[2] : y_lo[2];
    assign Y[1]   = v_hi ? y_hi[1] : y_lo[1];
    assign Y[0]   = v_hi ? y_hi[0] : y_lo[0];
